`timescale 1ns/1ns
`include "config.v"
module softmax_controller (
	input clk,
	input rst,
    input softmax_en,
    output is_stage2,
    output is_stage4
);
    reg [] cnt;
    

endmodule

